// The various set/read commands below have hard coded the relevant data.
// The data being set is in the final byte of the command. When reading,
// the last byte we send is irrelevant.

// Soft reset w5500
localparam SOFT_RESET_W5500 = 32'b00000000_00000000_00000100_10000000;

// Set PHY to 100 megabits / second, full duplex
localparam SET_PHY_MODE = 32'b00000000_00101110_00000100_11011000;


// Set/read our MAC address. 	SET: 	0x00 0x16 0x36 0xDE 0x58 0xF6
//										READ:	0x00 0x00 0x00 0xDE 0x58 0xF6
localparam SET_MAC_ADDRESS_BYTE_0  =  32'b00000000_00001001_00000100_00000000;
localparam READ_MAC_ADDRESS_BYTE_0 =  32'b00000000_00001001_00000000_00000000;
localparam SET_MAC_ADDRESS_BYTE_1  =  32'b00000000_00001010_00000100_00010110;
localparam READ_MAC_ADDRESS_BYTE_1 =  32'b00000000_00001010_00000000_00000000;
localparam SET_MAC_ADDRESS_BYTE_2  =  32'b00000000_00001011_00000100_00110110;
localparam READ_MAC_ADDRESS_BYTE_2 =  32'b00000000_00001011_00000000_00000000;
localparam SET_MAC_ADDRESS_BYTE_3  =  32'b00000000_00001100_00000100_11011110;
localparam READ_MAC_ADDRESS_BYTE_3 =  32'b00000000_00001100_00000000_11011110;
localparam SET_MAC_ADDRESS_BYTE_4  =  32'b00000000_00001101_00000100_01011000;
localparam READ_MAC_ADDRESS_BYTE_4 =  32'b00000000_00001101_00000000_01011000;
localparam SET_MAC_ADDRESS_BYTE_5  =  32'b00000000_00001110_00000100_11110110;
localparam READ_MAC_ADDRESS_BYTE_5 =  32'b00000000_00001110_00000000_11110110;

// Set/read our IP address. (192.168.0.12)
localparam SET_SOURCE_IP_ADDRESS_0  =  32'b00000000_00001111_00000100_11000000;
localparam READ_SOURCE_IP_ADDRESS_0 =  32'b00000000_00001111_00000000_00000000;
localparam SET_SOURCE_IP_ADDRESS_1  =  32'b00000000_00010000_00000100_10101000;
localparam READ_SOURCE_IP_ADDRESS_1 =  32'b00000000_00010000_00000000_00000000;
localparam SET_SOURCE_IP_ADDRESS_2  =  32'b00000000_00010001_00000100_00000000;
localparam READ_SOURCE_IP_ADDRESS_2 =  32'b00000000_00010001_00000000_00000000;
localparam SET_SOURCE_IP_ADDRESS_3  =  32'b00000000_00010010_00000100_00001100;
localparam READ_SOURCE_IP_ADDRESS_3 =  32'b00000000_00010010_00000000_00000000;

// Set/read out gateway address. (192.168.0.8)
localparam SET_GATEWAY_ADDRESS_0    = 32'b00000000_00000001_00000100_11000000;
localparam READ_GATEWAY_ADDRESS_0   = 32'b00000000_00000001_00000000_00000000;
localparam SET_GATEWAY_ADDRESS_1    = 32'b00000000_00000010_00000100_10101000;
localparam READ_GATEWAY_ADDRESS_1   = 32'b00000000_00000010_00000000_00000000;
localparam SET_GATEWAY_ADDRESS_2    = 32'b00000000_00000011_00000100_00000000;
localparam READ_GATEWAY_ADDRESS_2   = 32'b00000000_00000011_00000000_00000000;
localparam SET_GATEWAY_ADDRESS_3    = 32'b00000000_00000100_00000100_00001000;
localparam READ_GATEWAY_ADDRESS_3   = 32'b00000000_00000100_00000000_00000000;

// Set/read out subnet mask. (255.255.255.0)
localparam SET_SUBNET_MASK_0  = 32'b00000000_00000101_00000100_11111111;
localparam READ_SUBNET_MASK_0 = 32'b00000000_00000101_00000000_00000000;
localparam SET_SUBNET_MASK_1  = 32'b00000000_00000110_00000100_11111111;
localparam READ_SUBNET_MASK_1 = 32'b00000000_00000110_00000000_00000000;
localparam SET_SUBNET_MASK_2  = 32'b00000000_00000111_00000100_11111111;
localparam READ_SUBNET_MASK_2 = 32'b00000000_00000111_00000000_00000000;
localparam SET_SUBNET_MASK_3  = 32'b00000000_00001000_00000100_00000000;
localparam READ_SUBNET_MASK_3 = 32'b00000000_00001000_00000000_00000000;

// Set the socket mode to UDP with no blocking
localparam SET_SOCKET_0_MODE  = 32'b00000000_00000000_00001100_00000010;
localparam READ_SOCKET_0_MODE = 32'b00000000_00000000_00001000_00000010;

// Set the socket source port number to 5000. Requires two commands.
localparam SET_SOCKET_0_SRC_PORT_0 = 32'b00000000_00000100_00001100_00010011;
localparam SET_SOCKET_0_SRC_PORT_1 = 32'b00000000_00000101_00001100_10001000;

// Set socket 0's destination IP address (192.168.0.108) 
localparam SET_SOCKET_0_DST_IP_0 = 32'b00000000_00001100_00001100_11000000;
localparam SET_SOCKET_0_DST_IP_1 = 32'b00000000_00001101_00001100_10101000;
localparam SET_SOCKET_0_DST_IP_2 = 32'b00000000_00001110_00001100_00000000;
localparam SET_SOCKET_0_DST_IP_3 = 32'b00000000_00001111_00001100_01101100;

// Set socket 0's destination port to 5000. Requires two commands.
localparam SET_SOCKET_0_DST_PRT_0 = 32'b00000000_00010000_00001100_00010011;
localparam SET_SOCKET_0_DST_PRT_1 = 32'b00000000_00010001_00001100_10001000;

// Set socket 0's TX buffer size to 16kilobytes
localparam SET_SOCKET_0_TX_BFR_SZ = 32'b00000000_00011111_00001100_00010000;

localparam OPEN_SOCKET_0 = 32'b00000000_00000001_00001100_00000001;
localparam READ_SOCKET_0_STATE = 32'b00000000_00000011_00001000_00100010;


localparam SEND_PACKET_SOCKET_0 = 32'b00000000_00000001_00001100_00100000;
localparam READ_CHIP_VERSION       = 32'b00000000001110010000000000000000;